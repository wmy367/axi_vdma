/**********************************************
______________                ______________
______________ \  /\  /|\  /| ______________
______________  \/  \/ | \/ | ______________
descript:
    axi4 write read lock ,pend each other
author : Young
Version: VERA.0.0
creaded: 2016/8/29 下午3:29:24
madified:
***********************************************/
`timescale 1ns/1ps
module axi4_interconnect_wrap #(
    parameter AXI_DSIZE = 256
)(
    input          INTERCONNECT_ACLK    ,
    input          INTERCONNECT_ARESETN ,

    output         S00_AXI_ARESET_OUT_N ,
    output         S01_AXI_ARESET_OUT_N ,
    output         S02_AXI_ARESET_OUT_N ,
    output         S03_AXI_ARESET_OUT_N ,
    output         S04_AXI_ARESET_OUT_N ,
    output         S05_AXI_ARESET_OUT_N ,
    output         S06_AXI_ARESET_OUT_N ,
    output         S07_AXI_ARESET_OUT_N ,
    output         M00_AXI_ARESET_OUT_N ,
    axi_inf.slaver s00_inf  ,
    axi_inf.slaver s01_inf  ,
    axi_inf.slaver s02_inf  ,
    axi_inf.slaver s03_inf  ,
    axi_inf.slaver s04_inf  ,
    axi_inf.slaver s05_inf  ,
    axi_inf.slaver s06_inf  ,
    axi_inf.slaver s07_inf  ,
    axi_inf.master m00_inf
);

generate
if(AXI_DSIZE ==256)begin
AXI4_INFCNT AXI4_INFCNT_inst(
/*  input          */   .INTERCONNECT_ACLK               (INTERCONNECT_ACLK          ),
/*  input          */   .INTERCONNECT_ARESETN            (INTERCONNECT_ARESETN       ),
/*  output         */   .S00_AXI_ARESET_OUT_N            (S00_AXI_ARESET_OUT_N       ),
/*  input          */   .S00_AXI_ACLK                    (s00_inf.axi_aclk           ),
/*  input [0:0]    */   .S00_AXI_AWID                    (s00_inf.axi_awid           ),
/*  input [28:0]   */   .S00_AXI_AWADDR                  (s00_inf.axi_awaddr         ),
/*  input [7:0]    */   .S00_AXI_AWLEN                   (s00_inf.axi_awlen          ),
/*  input [2:0]    */   .S00_AXI_AWSIZE                  (s00_inf.axi_awsize         ),
/*  input [1:0]    */   .S00_AXI_AWBURST                 (s00_inf.axi_awburst        ),
/*  input          */   .S00_AXI_AWLOCK                  (s00_inf.axi_awlock         ),
/*  input [3:0]    */   .S00_AXI_AWCACHE                 (s00_inf.axi_awcache        ),
/*  input [2:0]    */   .S00_AXI_AWPROT                  (s00_inf.axi_awprot         ),
/*  input [3:0]    */   .S00_AXI_AWQOS                   (s00_inf.axi_awqos          ),
/*  input          */   .S00_AXI_AWVALID                 (s00_inf.axi_awvalid        ),
/*  output         */   .S00_AXI_AWREADY                 (s00_inf.axi_awready        ),
/*  input [255:0]  */   .S00_AXI_WDATA                   (s00_inf.axi_wdata          ),
/*  input [31:0]   */   .S00_AXI_WSTRB                   (s00_inf.axi_wstrb          ),
/*  input          */   .S00_AXI_WLAST                   (s00_inf.axi_wlast          ),
/*  input          */   .S00_AXI_WVALID                  (s00_inf.axi_wvalid         ),
/*  output         */   .S00_AXI_WREADY                  (s00_inf.axi_wready         ),
/*  output [0:0]   */   .S00_AXI_BID                     (s00_inf.axi_bid            ),
/*  output [1:0]   */   .S00_AXI_BRESP                   (s00_inf.axi_bresp          ),
/*  output         */   .S00_AXI_BVALID                  (s00_inf.axi_bvalid         ),
/*  input          */   .S00_AXI_BREADY                  (s00_inf.axi_bready         ),
/*  input [0:0]    */   .S00_AXI_ARID                    (s00_inf.axi_arid           ),
/*  input [28:0]   */   .S00_AXI_ARADDR                  (s00_inf.axi_araddr         ),
/*  input [7:0]    */   .S00_AXI_ARLEN                   (s00_inf.axi_arlen          ),
/*  input [2:0]    */   .S00_AXI_ARSIZE                  (s00_inf.axi_arsize         ),
/*  input [1:0]    */   .S00_AXI_ARBURST                 (s00_inf.axi_arburst        ),
/*  input          */   .S00_AXI_ARLOCK                  (s00_inf.axi_arlock         ),
/*  input [3:0]    */   .S00_AXI_ARCACHE                 (s00_inf.axi_arcache        ),
/*  input [2:0]    */   .S00_AXI_ARPROT                  (s00_inf.axi_arprot         ),
/*  input [3:0]    */   .S00_AXI_ARQOS                   (s00_inf.axi_arqos          ),
/*  input          */   .S00_AXI_ARVALID                 (s00_inf.axi_arvalid        ),
/*  output         */   .S00_AXI_ARREADY                 (s00_inf.axi_arready        ),
/*  output [0:0]   */   .S00_AXI_RID                     (s00_inf.axi_rid            ),
/*  output [255:0] */   .S00_AXI_RDATA                   (s00_inf.axi_rdata          ),
/*  output [1:0]   */   .S00_AXI_RRESP                   (s00_inf.axi_rresp          ),
/*  output         */   .S00_AXI_RLAST                   (s00_inf.axi_rlast          ),
/*  output         */   .S00_AXI_RVALID                  (s00_inf.axi_rvalid         ),
/*  input          */   .S00_AXI_RREADY                  (s00_inf.axi_rready         ),
/*  output S01_AXI_*/   .S01_AXI_ARESET_OUT_N            (S01_AXI_ARESET_OUT_N       ),
/*  input          */   .S01_AXI_ACLK                    (s01_inf.axi_aclk               ),
/*  input [0:0]    */   .S01_AXI_AWID                    (s01_inf.axi_awid               ),
/*  input [28:0]   */   .S01_AXI_AWADDR                  (s01_inf.axi_awaddr             ),
/*  input [7:0]    */   .S01_AXI_AWLEN                   (s01_inf.axi_awlen              ),
/*  input [2:0]    */   .S01_AXI_AWSIZE                  (s01_inf.axi_awsize             ),
/*  input [1:0]    */   .S01_AXI_AWBURST                 (s01_inf.axi_awburst            ),
/*  input          */   .S01_AXI_AWLOCK                  (s01_inf.axi_awlock             ),
/*  input [3:0]    */   .S01_AXI_AWCACHE                 (s01_inf.axi_awcache            ),
/*  input [2:0]    */   .S01_AXI_AWPROT                  (s01_inf.axi_awprot             ),
/*  input [3:0]    */   .S01_AXI_AWQOS                   (s01_inf.axi_awqos              ),
/*  input          */   .S01_AXI_AWVALID                 (s01_inf.axi_awvalid            ),
/*  output         */   .S01_AXI_AWREADY                 (s01_inf.axi_awready            ),
/*  input [255:0]  */   .S01_AXI_WDATA                   (s01_inf.axi_wdata              ),
/*  input [31:0]   */   .S01_AXI_WSTRB                   (s01_inf.axi_wstrb              ),
/*  input          */   .S01_AXI_WLAST                   (s01_inf.axi_wlast              ),
/*  input          */   .S01_AXI_WVALID                  (s01_inf.axi_wvalid             ),
/*  output         */   .S01_AXI_WREADY                  (s01_inf.axi_wready             ),
/*  output [0:0]   */   .S01_AXI_BID                     (s01_inf.axi_bid                ),
/*  output [1:0]   */   .S01_AXI_BRESP                   (s01_inf.axi_bresp              ),
/*  output         */   .S01_AXI_BVALID                  (s01_inf.axi_bvalid             ),
/*  input          */   .S01_AXI_BREADY                  (s01_inf.axi_bready             ),
/*  input [0:0]    */   .S01_AXI_ARID                    (s01_inf.axi_arid               ),
/*  input [28:0]   */   .S01_AXI_ARADDR                  (s01_inf.axi_araddr             ),
/*  input [7:0]    */   .S01_AXI_ARLEN                   (s01_inf.axi_arlen              ),
/*  input [2:0]    */   .S01_AXI_ARSIZE                  (s01_inf.axi_arsize             ),
/*  input [1:0]    */   .S01_AXI_ARBURST                 (s01_inf.axi_arburst            ),
/*  input          */   .S01_AXI_ARLOCK                  (s01_inf.axi_arlock             ),
/*  input [3:0]    */   .S01_AXI_ARCACHE                 (s01_inf.axi_arcache            ),
/*  input [2:0]    */   .S01_AXI_ARPROT                  (s01_inf.axi_arprot             ),
/*  input [3:0]    */   .S01_AXI_ARQOS                   (s01_inf.axi_arqos              ),
/*  input          */   .S01_AXI_ARVALID                 (s01_inf.axi_arvalid            ),
/*  output         */   .S01_AXI_ARREADY                 (s01_inf.axi_arready            ),
/*  output [0:0]   */   .S01_AXI_RID                     (s01_inf.axi_rid                ),
/*  output [255:0] */   .S01_AXI_RDATA                   (s01_inf.axi_rdata              ),
/*  output [1:0]   */   .S01_AXI_RRESP                   (s01_inf.axi_rresp              ),
/*  output         */   .S01_AXI_RLAST                   (s01_inf.axi_rlast              ),
/*  output         */   .S01_AXI_RVALID                  (s01_inf.axi_rvalid             ),
/*  input          */   .S01_AXI_RREADY                  (s01_inf.axi_rready             ),

/*  output         */   .S02_AXI_ARESET_OUT_N            (S02_AXI_ARESET_OUT_N       ),
/*  input          */   .S02_AXI_ACLK                    (s02_inf.axi_aclk           ),
/*  input [0:0]    */   .S02_AXI_AWID                    (s02_inf.axi_awid           ),
/*  input [28:0]   */   .S02_AXI_AWADDR                  (s02_inf.axi_awaddr         ),
/*  input [7:0]    */   .S02_AXI_AWLEN                   (s02_inf.axi_awlen          ),
/*  input [2:0]    */   .S02_AXI_AWSIZE                  (s02_inf.axi_awsize         ),
/*  input [1:0]    */   .S02_AXI_AWBURST                 (s02_inf.axi_awburst        ),
/*  input          */   .S02_AXI_AWLOCK                  (s02_inf.axi_awlock         ),
/*  input [3:0]    */   .S02_AXI_AWCACHE                 (s02_inf.axi_awcache        ),
/*  input [2:0]    */   .S02_AXI_AWPROT                  (s02_inf.axi_awprot         ),
/*  input [3:0]    */   .S02_AXI_AWQOS                   (s02_inf.axi_awqos          ),
/*  input          */   .S02_AXI_AWVALID                 (s02_inf.axi_awvalid        ),
/*  output         */   .S02_AXI_AWREADY                 (s02_inf.axi_awready        ),
/*  input [255:0]  */   .S02_AXI_WDATA                   (s02_inf.axi_wdata          ),
/*  input [31:0]   */   .S02_AXI_WSTRB                   (s02_inf.axi_wstrb          ),
/*  input          */   .S02_AXI_WLAST                   (s02_inf.axi_wlast          ),
/*  input          */   .S02_AXI_WVALID                  (s02_inf.axi_wvalid         ),
/*  output         */   .S02_AXI_WREADY                  (s02_inf.axi_wready         ),
/*  output [0:0]   */   .S02_AXI_BID                     (s02_inf.axi_bid            ),
/*  output [1:0]   */   .S02_AXI_BRESP                   (s02_inf.axi_bresp          ),
/*  output         */   .S02_AXI_BVALID                  (s02_inf.axi_bvalid         ),
/*  input          */   .S02_AXI_BREADY                  (s02_inf.axi_bready         ),
/*  input [0:0]    */   .S02_AXI_ARID                    (s02_inf.axi_arid           ),
/*  input [28:0]   */   .S02_AXI_ARADDR                  (s02_inf.axi_araddr         ),
/*  input [7:0]    */   .S02_AXI_ARLEN                   (s02_inf.axi_arlen          ),
/*  input [2:0]    */   .S02_AXI_ARSIZE                  (s02_inf.axi_arsize         ),
/*  input [1:0]    */   .S02_AXI_ARBURST                 (s02_inf.axi_arburst        ),
/*  input          */   .S02_AXI_ARLOCK                  (s02_inf.axi_arlock         ),
/*  input [3:0]    */   .S02_AXI_ARCACHE                 (s02_inf.axi_arcache        ),
/*  input [2:0]    */   .S02_AXI_ARPROT                  (s02_inf.axi_arprot         ),
/*  input [3:0]    */   .S02_AXI_ARQOS                   (s02_inf.axi_arqos          ),
/*  input          */   .S02_AXI_ARVALID                 (s02_inf.axi_arvalid        ),
/*  output         */   .S02_AXI_ARREADY                 (s02_inf.axi_arready        ),
/*  output [0:0]   */   .S02_AXI_RID                     (s02_inf.axi_rid            ),
/*  output [255:0] */   .S02_AXI_RDATA                   (s02_inf.axi_rdata          ),
/*  output [1:0]   */   .S02_AXI_RRESP                   (s02_inf.axi_rresp          ),
/*  output         */   .S02_AXI_RLAST                   (s02_inf.axi_rlast          ),
/*  output         */   .S02_AXI_RVALID                  (s02_inf.axi_rvalid         ),
/*  input          */   .S02_AXI_RREADY                  (s02_inf.axi_rready         ),
/*  output S01_AXI_*/   .S03_AXI_ARESET_OUT_N            (S03_AXI_ARESET_OUT_N       ),
/*  input          */   .S03_AXI_ACLK                    (s03_inf.axi_aclk               ),
/*  input [0:0]    */   .S03_AXI_AWID                    (s03_inf.axi_awid               ),
/*  input [28:0]   */   .S03_AXI_AWADDR                  (s03_inf.axi_awaddr             ),
/*  input [7:0]    */   .S03_AXI_AWLEN                   (s03_inf.axi_awlen              ),
/*  input [2:0]    */   .S03_AXI_AWSIZE                  (s03_inf.axi_awsize             ),
/*  input [1:0]    */   .S03_AXI_AWBURST                 (s03_inf.axi_awburst            ),
/*  input          */   .S03_AXI_AWLOCK                  (s03_inf.axi_awlock             ),
/*  input [3:0]    */   .S03_AXI_AWCACHE                 (s03_inf.axi_awcache            ),
/*  input [2:0]    */   .S03_AXI_AWPROT                  (s03_inf.axi_awprot             ),
/*  input [3:0]    */   .S03_AXI_AWQOS                   (s03_inf.axi_awqos              ),
/*  input          */   .S03_AXI_AWVALID                 (s03_inf.axi_awvalid            ),
/*  output         */   .S03_AXI_AWREADY                 (s03_inf.axi_awready            ),
/*  input [255:0]  */   .S03_AXI_WDATA                   (s03_inf.axi_wdata              ),
/*  input [31:0]   */   .S03_AXI_WSTRB                   (s03_inf.axi_wstrb              ),
/*  input          */   .S03_AXI_WLAST                   (s03_inf.axi_wlast              ),
/*  input          */   .S03_AXI_WVALID                  (s03_inf.axi_wvalid             ),
/*  output         */   .S03_AXI_WREADY                  (s03_inf.axi_wready             ),
/*  output [0:0]   */   .S03_AXI_BID                     (s03_inf.axi_bid                ),
/*  output [1:0]   */   .S03_AXI_BRESP                   (s03_inf.axi_bresp              ),
/*  output         */   .S03_AXI_BVALID                  (s03_inf.axi_bvalid             ),
/*  input          */   .S03_AXI_BREADY                  (s03_inf.axi_bready             ),
/*  input [0:0]    */   .S03_AXI_ARID                    (s03_inf.axi_arid               ),
/*  input [28:0]   */   .S03_AXI_ARADDR                  (s03_inf.axi_araddr             ),
/*  input [7:0]    */   .S03_AXI_ARLEN                   (s03_inf.axi_arlen              ),
/*  input [2:0]    */   .S03_AXI_ARSIZE                  (s03_inf.axi_arsize             ),
/*  input [1:0]    */   .S03_AXI_ARBURST                 (s03_inf.axi_arburst            ),
/*  input          */   .S03_AXI_ARLOCK                  (s03_inf.axi_arlock             ),
/*  input [3:0]    */   .S03_AXI_ARCACHE                 (s03_inf.axi_arcache            ),
/*  input [2:0]    */   .S03_AXI_ARPROT                  (s03_inf.axi_arprot             ),
/*  input [3:0]    */   .S03_AXI_ARQOS                   (s03_inf.axi_arqos              ),
/*  input          */   .S03_AXI_ARVALID                 (s03_inf.axi_arvalid            ),
/*  output         */   .S03_AXI_ARREADY                 (s03_inf.axi_arready            ),
/*  output [0:0]   */   .S03_AXI_RID                     (s03_inf.axi_rid                ),
/*  output [255:0] */   .S03_AXI_RDATA                   (s03_inf.axi_rdata              ),
/*  output [1:0]   */   .S03_AXI_RRESP                   (s03_inf.axi_rresp              ),
/*  output         */   .S03_AXI_RLAST                   (s03_inf.axi_rlast              ),
/*  output         */   .S03_AXI_RVALID                  (s03_inf.axi_rvalid             ),
/*  input          */   .S03_AXI_RREADY                  (s03_inf.axi_rready             ),

/*  output         */   .S04_AXI_ARESET_OUT_N            (S04_AXI_ARESET_OUT_N       ),
/*  input          */   .S04_AXI_ACLK                    (s04_inf.axi_aclk           ),
/*  input [0:0]    */   .S04_AXI_AWID                    (s04_inf.axi_awid           ),
/*  input [28:0]   */   .S04_AXI_AWADDR                  (s04_inf.axi_awaddr         ),
/*  input [7:0]    */   .S04_AXI_AWLEN                   (s04_inf.axi_awlen          ),
/*  input [2:0]    */   .S04_AXI_AWSIZE                  (s04_inf.axi_awsize         ),
/*  input [1:0]    */   .S04_AXI_AWBURST                 (s04_inf.axi_awburst        ),
/*  input          */   .S04_AXI_AWLOCK                  (s04_inf.axi_awlock         ),
/*  input [3:0]    */   .S04_AXI_AWCACHE                 (s04_inf.axi_awcache        ),
/*  input [2:0]    */   .S04_AXI_AWPROT                  (s04_inf.axi_awprot         ),
/*  input [3:0]    */   .S04_AXI_AWQOS                   (s04_inf.axi_awqos          ),
/*  input          */   .S04_AXI_AWVALID                 (s04_inf.axi_awvalid        ),
/*  output         */   .S04_AXI_AWREADY                 (s04_inf.axi_awready        ),
/*  input [255:0]  */   .S04_AXI_WDATA                   (s04_inf.axi_wdata          ),
/*  input [31:0]   */   .S04_AXI_WSTRB                   (s04_inf.axi_wstrb          ),
/*  input          */   .S04_AXI_WLAST                   (s04_inf.axi_wlast          ),
/*  input          */   .S04_AXI_WVALID                  (s04_inf.axi_wvalid         ),
/*  output         */   .S04_AXI_WREADY                  (s04_inf.axi_wready         ),
/*  output [0:0]   */   .S04_AXI_BID                     (s04_inf.axi_bid            ),
/*  output [1:0]   */   .S04_AXI_BRESP                   (s04_inf.axi_bresp          ),
/*  output         */   .S04_AXI_BVALID                  (s04_inf.axi_bvalid         ),
/*  input          */   .S04_AXI_BREADY                  (s04_inf.axi_bready         ),
/*  input [0:0]    */   .S04_AXI_ARID                    (s04_inf.axi_arid           ),
/*  input [28:0]   */   .S04_AXI_ARADDR                  (s04_inf.axi_araddr         ),
/*  input [7:0]    */   .S04_AXI_ARLEN                   (s04_inf.axi_arlen          ),
/*  input [2:0]    */   .S04_AXI_ARSIZE                  (s04_inf.axi_arsize         ),
/*  input [1:0]    */   .S04_AXI_ARBURST                 (s04_inf.axi_arburst        ),
/*  input          */   .S04_AXI_ARLOCK                  (s04_inf.axi_arlock         ),
/*  input [3:0]    */   .S04_AXI_ARCACHE                 (s04_inf.axi_arcache        ),
/*  input [2:0]    */   .S04_AXI_ARPROT                  (s04_inf.axi_arprot         ),
/*  input [3:0]    */   .S04_AXI_ARQOS                   (s04_inf.axi_arqos          ),
/*  input          */   .S04_AXI_ARVALID                 (s04_inf.axi_arvalid        ),
/*  output         */   .S04_AXI_ARREADY                 (s04_inf.axi_arready        ),
/*  output [0:0]   */   .S04_AXI_RID                     (s04_inf.axi_rid            ),
/*  output [255:0] */   .S04_AXI_RDATA                   (s04_inf.axi_rdata          ),
/*  output [1:0]   */   .S04_AXI_RRESP                   (s04_inf.axi_rresp          ),
/*  output         */   .S04_AXI_RLAST                   (s04_inf.axi_rlast          ),
/*  output         */   .S04_AXI_RVALID                  (s04_inf.axi_rvalid         ),
/*  input          */   .S04_AXI_RREADY                  (s04_inf.axi_rready         ),
/*  output S01_AXI_*/   .S05_AXI_ARESET_OUT_N            (S05_AXI_ARESET_OUT_N       ),
/*  input          */   .S05_AXI_ACLK                    (s05_inf.axi_aclk               ),
/*  input [0:0]    */   .S05_AXI_AWID                    (s05_inf.axi_awid               ),
/*  input [28:0]   */   .S05_AXI_AWADDR                  (s05_inf.axi_awaddr             ),
/*  input [7:0]    */   .S05_AXI_AWLEN                   (s05_inf.axi_awlen              ),
/*  input [2:0]    */   .S05_AXI_AWSIZE                  (s05_inf.axi_awsize             ),
/*  input [1:0]    */   .S05_AXI_AWBURST                 (s05_inf.axi_awburst            ),
/*  input          */   .S05_AXI_AWLOCK                  (s05_inf.axi_awlock             ),
/*  input [3:0]    */   .S05_AXI_AWCACHE                 (s05_inf.axi_awcache            ),
/*  input [2:0]    */   .S05_AXI_AWPROT                  (s05_inf.axi_awprot             ),
/*  input [3:0]    */   .S05_AXI_AWQOS                   (s05_inf.axi_awqos              ),
/*  input          */   .S05_AXI_AWVALID                 (s05_inf.axi_awvalid            ),
/*  output         */   .S05_AXI_AWREADY                 (s05_inf.axi_awready            ),
/*  input [255:0]  */   .S05_AXI_WDATA                   (s05_inf.axi_wdata              ),
/*  input [31:0]   */   .S05_AXI_WSTRB                   (s05_inf.axi_wstrb              ),
/*  input          */   .S05_AXI_WLAST                   (s05_inf.axi_wlast              ),
/*  input          */   .S05_AXI_WVALID                  (s05_inf.axi_wvalid             ),
/*  output         */   .S05_AXI_WREADY                  (s05_inf.axi_wready             ),
/*  output [0:0]   */   .S05_AXI_BID                     (s05_inf.axi_bid                ),
/*  output [1:0]   */   .S05_AXI_BRESP                   (s05_inf.axi_bresp              ),
/*  output         */   .S05_AXI_BVALID                  (s05_inf.axi_bvalid             ),
/*  input          */   .S05_AXI_BREADY                  (s05_inf.axi_bready             ),
/*  input [0:0]    */   .S05_AXI_ARID                    (s05_inf.axi_arid               ),
/*  input [28:0]   */   .S05_AXI_ARADDR                  (s05_inf.axi_araddr             ),
/*  input [7:0]    */   .S05_AXI_ARLEN                   (s05_inf.axi_arlen              ),
/*  input [2:0]    */   .S05_AXI_ARSIZE                  (s05_inf.axi_arsize             ),
/*  input [1:0]    */   .S05_AXI_ARBURST                 (s05_inf.axi_arburst            ),
/*  input          */   .S05_AXI_ARLOCK                  (s05_inf.axi_arlock             ),
/*  input [3:0]    */   .S05_AXI_ARCACHE                 (s05_inf.axi_arcache            ),
/*  input [2:0]    */   .S05_AXI_ARPROT                  (s05_inf.axi_arprot             ),
/*  input [3:0]    */   .S05_AXI_ARQOS                   (s05_inf.axi_arqos              ),
/*  input          */   .S05_AXI_ARVALID                 (s05_inf.axi_arvalid            ),
/*  output         */   .S05_AXI_ARREADY                 (s05_inf.axi_arready            ),
/*  output [0:0]   */   .S05_AXI_RID                     (s05_inf.axi_rid                ),
/*  output [255:0] */   .S05_AXI_RDATA                   (s05_inf.axi_rdata              ),
/*  output [1:0]   */   .S05_AXI_RRESP                   (s05_inf.axi_rresp              ),
/*  output         */   .S05_AXI_RLAST                   (s05_inf.axi_rlast              ),
/*  output         */   .S05_AXI_RVALID                  (s05_inf.axi_rvalid             ),
/*  input          */   .S05_AXI_RREADY                  (s05_inf.axi_rready             ),

/*  output         */   .S06_AXI_ARESET_OUT_N            (S06_AXI_ARESET_OUT_N       ),
/*  input          */   .S06_AXI_ACLK                    (s06_inf.axi_aclk           ),
/*  input [0:0]    */   .S06_AXI_AWID                    (s06_inf.axi_awid           ),
/*  input [28:0]   */   .S06_AXI_AWADDR                  (s06_inf.axi_awaddr         ),
/*  input [7:0]    */   .S06_AXI_AWLEN                   (s06_inf.axi_awlen          ),
/*  input [2:0]    */   .S06_AXI_AWSIZE                  (s06_inf.axi_awsize         ),
/*  input [1:0]    */   .S06_AXI_AWBURST                 (s06_inf.axi_awburst        ),
/*  input          */   .S06_AXI_AWLOCK                  (s06_inf.axi_awlock         ),
/*  input [3:0]    */   .S06_AXI_AWCACHE                 (s06_inf.axi_awcache        ),
/*  input [2:0]    */   .S06_AXI_AWPROT                  (s06_inf.axi_awprot         ),
/*  input [3:0]    */   .S06_AXI_AWQOS                   (s06_inf.axi_awqos          ),
/*  input          */   .S06_AXI_AWVALID                 (s06_inf.axi_awvalid        ),
/*  output         */   .S06_AXI_AWREADY                 (s06_inf.axi_awready        ),
/*  input [255:0]  */   .S06_AXI_WDATA                   (s06_inf.axi_wdata          ),
/*  input [31:0]   */   .S06_AXI_WSTRB                   (s06_inf.axi_wstrb          ),
/*  input          */   .S06_AXI_WLAST                   (s06_inf.axi_wlast          ),
/*  input          */   .S06_AXI_WVALID                  (s06_inf.axi_wvalid         ),
/*  output         */   .S06_AXI_WREADY                  (s06_inf.axi_wready         ),
/*  output [0:0]   */   .S06_AXI_BID                     (s06_inf.axi_bid            ),
/*  output [1:0]   */   .S06_AXI_BRESP                   (s06_inf.axi_bresp          ),
/*  output         */   .S06_AXI_BVALID                  (s06_inf.axi_bvalid         ),
/*  input          */   .S06_AXI_BREADY                  (s06_inf.axi_bready         ),
/*  input [0:0]    */   .S06_AXI_ARID                    (s06_inf.axi_arid           ),
/*  input [28:0]   */   .S06_AXI_ARADDR                  (s06_inf.axi_araddr         ),
/*  input [7:0]    */   .S06_AXI_ARLEN                   (s06_inf.axi_arlen          ),
/*  input [2:0]    */   .S06_AXI_ARSIZE                  (s06_inf.axi_arsize         ),
/*  input [1:0]    */   .S06_AXI_ARBURST                 (s06_inf.axi_arburst        ),
/*  input          */   .S06_AXI_ARLOCK                  (s06_inf.axi_arlock         ),
/*  input [3:0]    */   .S06_AXI_ARCACHE                 (s06_inf.axi_arcache        ),
/*  input [2:0]    */   .S06_AXI_ARPROT                  (s06_inf.axi_arprot         ),
/*  input [3:0]    */   .S06_AXI_ARQOS                   (s06_inf.axi_arqos          ),
/*  input          */   .S06_AXI_ARVALID                 (s06_inf.axi_arvalid        ),
/*  output         */   .S06_AXI_ARREADY                 (s06_inf.axi_arready        ),
/*  output [0:0]   */   .S06_AXI_RID                     (s06_inf.axi_rid            ),
/*  output [255:0] */   .S06_AXI_RDATA                   (s06_inf.axi_rdata          ),
/*  output [1:0]   */   .S06_AXI_RRESP                   (s06_inf.axi_rresp          ),
/*  output         */   .S06_AXI_RLAST                   (s06_inf.axi_rlast          ),
/*  output         */   .S06_AXI_RVALID                  (s06_inf.axi_rvalid         ),
/*  input          */   .S06_AXI_RREADY                  (s06_inf.axi_rready         ),
/*  output S01_AXI_*/   .S07_AXI_ARESET_OUT_N            (S07_AXI_ARESET_OUT_N       ),
/*  input          */   .S07_AXI_ACLK                    (s07_inf.axi_aclk               ),
/*  input [0:0]    */   .S07_AXI_AWID                    (s07_inf.axi_awid               ),
/*  input [28:0]   */   .S07_AXI_AWADDR                  (s07_inf.axi_awaddr             ),
/*  input [7:0]    */   .S07_AXI_AWLEN                   (s07_inf.axi_awlen              ),
/*  input [2:0]    */   .S07_AXI_AWSIZE                  (s07_inf.axi_awsize             ),
/*  input [1:0]    */   .S07_AXI_AWBURST                 (s07_inf.axi_awburst            ),
/*  input          */   .S07_AXI_AWLOCK                  (s07_inf.axi_awlock             ),
/*  input [3:0]    */   .S07_AXI_AWCACHE                 (s07_inf.axi_awcache            ),
/*  input [2:0]    */   .S07_AXI_AWPROT                  (s07_inf.axi_awprot             ),
/*  input [3:0]    */   .S07_AXI_AWQOS                   (s07_inf.axi_awqos              ),
/*  input          */   .S07_AXI_AWVALID                 (s07_inf.axi_awvalid            ),
/*  output         */   .S07_AXI_AWREADY                 (s07_inf.axi_awready            ),
/*  input [255:0]  */   .S07_AXI_WDATA                   (s07_inf.axi_wdata              ),
/*  input [31:0]   */   .S07_AXI_WSTRB                   (s07_inf.axi_wstrb              ),
/*  input          */   .S07_AXI_WLAST                   (s07_inf.axi_wlast              ),
/*  input          */   .S07_AXI_WVALID                  (s07_inf.axi_wvalid             ),
/*  output         */   .S07_AXI_WREADY                  (s07_inf.axi_wready             ),
/*  output [0:0]   */   .S07_AXI_BID                     (s07_inf.axi_bid                ),
/*  output [1:0]   */   .S07_AXI_BRESP                   (s07_inf.axi_bresp              ),
/*  output         */   .S07_AXI_BVALID                  (s07_inf.axi_bvalid             ),
/*  input          */   .S07_AXI_BREADY                  (s07_inf.axi_bready             ),
/*  input [0:0]    */   .S07_AXI_ARID                    (s07_inf.axi_arid               ),
/*  input [28:0]   */   .S07_AXI_ARADDR                  (s07_inf.axi_araddr             ),
/*  input [7:0]    */   .S07_AXI_ARLEN                   (s07_inf.axi_arlen              ),
/*  input [2:0]    */   .S07_AXI_ARSIZE                  (s07_inf.axi_arsize             ),
/*  input [1:0]    */   .S07_AXI_ARBURST                 (s07_inf.axi_arburst            ),
/*  input          */   .S07_AXI_ARLOCK                  (s07_inf.axi_arlock             ),
/*  input [3:0]    */   .S07_AXI_ARCACHE                 (s07_inf.axi_arcache            ),
/*  input [2:0]    */   .S07_AXI_ARPROT                  (s07_inf.axi_arprot             ),
/*  input [3:0]    */   .S07_AXI_ARQOS                   (s07_inf.axi_arqos              ),
/*  input          */   .S07_AXI_ARVALID                 (s07_inf.axi_arvalid            ),
/*  output         */   .S07_AXI_ARREADY                 (s07_inf.axi_arready            ),
/*  output [0:0]   */   .S07_AXI_RID                     (s07_inf.axi_rid                ),
/*  output [255:0] */   .S07_AXI_RDATA                   (s07_inf.axi_rdata              ),
/*  output [1:0]   */   .S07_AXI_RRESP                   (s07_inf.axi_rresp              ),
/*  output         */   .S07_AXI_RLAST                   (s07_inf.axi_rlast              ),
/*  output         */   .S07_AXI_RVALID                  (s07_inf.axi_rvalid             ),
/*  input          */   .S07_AXI_RREADY                  (s07_inf.axi_rready             ),


/*  output         */   .M00_AXI_ARESET_OUT_N            (M00_AXI_ARESET_OUT_N           ),
/*  input          */   .M00_AXI_ACLK                    (m00_inf.axi_aclk               ),
/*  output [3:0]   */   .M00_AXI_AWID                    (m00_inf.axi_awid               ),
/*  output [28:0]  */   .M00_AXI_AWADDR                  (m00_inf.axi_awaddr             ),
/*  output [7:0]   */   .M00_AXI_AWLEN                   (m00_inf.axi_awlen              ),
/*  output [2:0]   */   .M00_AXI_AWSIZE                  (m00_inf.axi_awsize             ),
/*  output [1:0]   */   .M00_AXI_AWBURST                 (m00_inf.axi_awburst            ),
/*  output         */   .M00_AXI_AWLOCK                  (m00_inf.axi_awlock             ),
/*  output [3:0]   */   .M00_AXI_AWCACHE                 (m00_inf.axi_awcache            ),
/*  output [2:0]   */   .M00_AXI_AWPROT                  (m00_inf.axi_awprot             ),
/*  output [3:0]   */   .M00_AXI_AWQOS                   (m00_inf.axi_awqos              ),
/*  output         */   .M00_AXI_AWVALID                 (m00_inf.axi_awvalid            ),
/*  input          */   .M00_AXI_AWREADY                 (m00_inf.axi_awready            ),
/*  output [255:0] */   .M00_AXI_WDATA                   (m00_inf.axi_wdata              ),
/*  output [31:0]  */   .M00_AXI_WSTRB                   (m00_inf.axi_wstrb              ),
/*  output         */   .M00_AXI_WLAST                   (m00_inf.axi_wlast              ),
/*  output         */   .M00_AXI_WVALID                  (m00_inf.axi_wvalid             ),
/*  input          */   .M00_AXI_WREADY                  (m00_inf.axi_wready             ),
/*  input [3:0]    */   .M00_AXI_BID                     (m00_inf.axi_bid                ),
/*  input [1:0]    */   .M00_AXI_BRESP                   (m00_inf.axi_bresp              ),
/*  input          */   .M00_AXI_BVALID                  (m00_inf.axi_bvalid             ),
/*  output         */   .M00_AXI_BREADY                  (m00_inf.axi_bready             ),
/*  output [3:0]   */   .M00_AXI_ARID                    (m00_inf.axi_arid               ),
/*  output [28:0]  */   .M00_AXI_ARADDR                  (m00_inf.axi_araddr             ),
/*  output [7:0]   */   .M00_AXI_ARLEN                   (m00_inf.axi_arlen              ),
/*  output [2:0]   */   .M00_AXI_ARSIZE                  (m00_inf.axi_arsize             ),
/*  output [1:0]   */   .M00_AXI_ARBURST                 (m00_inf.axi_arburst            ),
/*  output         */   .M00_AXI_ARLOCK                  (m00_inf.axi_arlock             ),
/*  output [3:0]   */   .M00_AXI_ARCACHE                 (m00_inf.axi_arcache            ),
/*  output [2:0]   */   .M00_AXI_ARPROT                  (m00_inf.axi_arprot             ),
/*  output [3:0]   */   .M00_AXI_ARQOS                   (m00_inf.axi_arqos              ),
/*  output         */   .M00_AXI_ARVALID                 (m00_inf.axi_arvalid            ),
/*  input          */   .M00_AXI_ARREADY                 (m00_inf.axi_arready            ),
/*  input [3:0]    */   .M00_AXI_RID                     (m00_inf.axi_rid                ),
/*  input [255:0]  */   .M00_AXI_RDATA                   (m00_inf.axi_rdata              ),
/*  input [1:0]    */   .M00_AXI_RRESP                   (m00_inf.axi_rresp              ),
/*  input          */   .M00_AXI_RLAST                   (m00_inf.axi_rlast              ),
/*  input          */   .M00_AXI_RVALID                  (m00_inf.axi_rvalid             ),
/*  output         */   .M00_AXI_RREADY                  (m00_inf.axi_rready             )
);
end else if(AXI_DSIZE == 512)begin
AXI4_INFCNT_512 AXI4_INFCNT_inst(
/*  input          */   .INTERCONNECT_ACLK               (INTERCONNECT_ACLK          ),
/*  input          */   .INTERCONNECT_ARESETN            (INTERCONNECT_ARESETN       ),
/*  output         */   .S00_AXI_ARESET_OUT_N            (S00_AXI_ARESET_OUT_N       ),
/*  input          */   .S00_AXI_ACLK                    (s00_inf.axi_aclk           ),
/*  input [0:0]    */   .S00_AXI_AWID                    (s00_inf.axi_awid           ),
/*  input [28:0]   */   .S00_AXI_AWADDR                  (s00_inf.axi_awaddr         ),
/*  input [7:0]    */   .S00_AXI_AWLEN                   (s00_inf.axi_awlen          ),
/*  input [2:0]    */   .S00_AXI_AWSIZE                  (s00_inf.axi_awsize         ),
/*  input [1:0]    */   .S00_AXI_AWBURST                 (s00_inf.axi_awburst        ),
/*  input          */   .S00_AXI_AWLOCK                  (s00_inf.axi_awlock         ),
/*  input [3:0]    */   .S00_AXI_AWCACHE                 (s00_inf.axi_awcache        ),
/*  input [2:0]    */   .S00_AXI_AWPROT                  (s00_inf.axi_awprot         ),
/*  input [3:0]    */   .S00_AXI_AWQOS                   (s00_inf.axi_awqos          ),
/*  input          */   .S00_AXI_AWVALID                 (s00_inf.axi_awvalid        ),
/*  output         */   .S00_AXI_AWREADY                 (s00_inf.axi_awready        ),
/*  input [511:0]  */   .S00_AXI_WDATA                   (s00_inf.axi_wdata          ),
/*  input [63:0]   */   .S00_AXI_WSTRB                   (s00_inf.axi_wstrb          ),
/*  input          */   .S00_AXI_WLAST                   (s00_inf.axi_wlast          ),
/*  input          */   .S00_AXI_WVALID                  (s00_inf.axi_wvalid         ),
/*  output         */   .S00_AXI_WREADY                  (s00_inf.axi_wready         ),
/*  output [0:0]   */   .S00_AXI_BID                     (s00_inf.axi_bid            ),
/*  output [1:0]   */   .S00_AXI_BRESP                   (s00_inf.axi_bresp          ),
/*  output         */   .S00_AXI_BVALID                  (s00_inf.axi_bvalid         ),
/*  input          */   .S00_AXI_BREADY                  (s00_inf.axi_bready         ),
/*  input [0:0]    */   .S00_AXI_ARID                    (s00_inf.axi_arid           ),
/*  input [28:0]   */   .S00_AXI_ARADDR                  (s00_inf.axi_araddr         ),
/*  input [7:0]    */   .S00_AXI_ARLEN                   (s00_inf.axi_arlen          ),
/*  input [2:0]    */   .S00_AXI_ARSIZE                  (s00_inf.axi_arsize         ),
/*  input [1:0]    */   .S00_AXI_ARBURST                 (s00_inf.axi_arburst        ),
/*  input          */   .S00_AXI_ARLOCK                  (s00_inf.axi_arlock         ),
/*  input [3:0]    */   .S00_AXI_ARCACHE                 (s00_inf.axi_arcache        ),
/*  input [2:0]    */   .S00_AXI_ARPROT                  (s00_inf.axi_arprot         ),
/*  input [3:0]    */   .S00_AXI_ARQOS                   (s00_inf.axi_arqos          ),
/*  input          */   .S00_AXI_ARVALID                 (s00_inf.axi_arvalid        ),
/*  output         */   .S00_AXI_ARREADY                 (s00_inf.axi_arready        ),
/*  output [0:0]   */   .S00_AXI_RID                     (s00_inf.axi_rid            ),
/*  output [511:0] */   .S00_AXI_RDATA                   (s00_inf.axi_rdata          ),
/*  output [1:0]   */   .S00_AXI_RRESP                   (s00_inf.axi_rresp          ),
/*  output         */   .S00_AXI_RLAST                   (s00_inf.axi_rlast          ),
/*  output         */   .S00_AXI_RVALID                  (s00_inf.axi_rvalid         ),
/*  input          */   .S00_AXI_RREADY                  (s00_inf.axi_rready         ),
/*  output S01_AXI_*/   .S01_AXI_ARESET_OUT_N            (S01_AXI_ARESET_OUT_N       ),
/*  input          */   .S01_AXI_ACLK                    (s01_inf.axi_aclk               ),
/*  input [0:0]    */   .S01_AXI_AWID                    (s01_inf.axi_awid               ),
/*  input [28:0]   */   .S01_AXI_AWADDR                  (s01_inf.axi_awaddr             ),
/*  input [7:0]    */   .S01_AXI_AWLEN                   (s01_inf.axi_awlen              ),
/*  input [2:0]    */   .S01_AXI_AWSIZE                  (s01_inf.axi_awsize             ),
/*  input [1:0]    */   .S01_AXI_AWBURST                 (s01_inf.axi_awburst            ),
/*  input          */   .S01_AXI_AWLOCK                  (s01_inf.axi_awlock             ),
/*  input [3:0]    */   .S01_AXI_AWCACHE                 (s01_inf.axi_awcache            ),
/*  input [2:0]    */   .S01_AXI_AWPROT                  (s01_inf.axi_awprot             ),
/*  input [3:0]    */   .S01_AXI_AWQOS                   (s01_inf.axi_awqos              ),
/*  input          */   .S01_AXI_AWVALID                 (s01_inf.axi_awvalid            ),
/*  output         */   .S01_AXI_AWREADY                 (s01_inf.axi_awready            ),
/*  input [511:0]  */   .S01_AXI_WDATA                   (s01_inf.axi_wdata              ),
/*  input [63:0]   */   .S01_AXI_WSTRB                   (s01_inf.axi_wstrb              ),
/*  input          */   .S01_AXI_WLAST                   (s01_inf.axi_wlast              ),
/*  input          */   .S01_AXI_WVALID                  (s01_inf.axi_wvalid             ),
/*  output         */   .S01_AXI_WREADY                  (s01_inf.axi_wready             ),
/*  output [0:0]   */   .S01_AXI_BID                     (s01_inf.axi_bid                ),
/*  output [1:0]   */   .S01_AXI_BRESP                   (s01_inf.axi_bresp              ),
/*  output         */   .S01_AXI_BVALID                  (s01_inf.axi_bvalid             ),
/*  input          */   .S01_AXI_BREADY                  (s01_inf.axi_bready             ),
/*  input [0:0]    */   .S01_AXI_ARID                    (s01_inf.axi_arid               ),
/*  input [28:0]   */   .S01_AXI_ARADDR                  (s01_inf.axi_araddr             ),
/*  input [7:0]    */   .S01_AXI_ARLEN                   (s01_inf.axi_arlen              ),
/*  input [2:0]    */   .S01_AXI_ARSIZE                  (s01_inf.axi_arsize             ),
/*  input [1:0]    */   .S01_AXI_ARBURST                 (s01_inf.axi_arburst            ),
/*  input          */   .S01_AXI_ARLOCK                  (s01_inf.axi_arlock             ),
/*  input [3:0]    */   .S01_AXI_ARCACHE                 (s01_inf.axi_arcache            ),
/*  input [2:0]    */   .S01_AXI_ARPROT                  (s01_inf.axi_arprot             ),
/*  input [3:0]    */   .S01_AXI_ARQOS                   (s01_inf.axi_arqos              ),
/*  input          */   .S01_AXI_ARVALID                 (s01_inf.axi_arvalid            ),
/*  output         */   .S01_AXI_ARREADY                 (s01_inf.axi_arready            ),
/*  output [0:0]   */   .S01_AXI_RID                     (s01_inf.axi_rid                ),
/*  output [511:0] */   .S01_AXI_RDATA                   (s01_inf.axi_rdata              ),
/*  output [1:0]   */   .S01_AXI_RRESP                   (s01_inf.axi_rresp              ),
/*  output         */   .S01_AXI_RLAST                   (s01_inf.axi_rlast              ),
/*  output         */   .S01_AXI_RVALID                  (s01_inf.axi_rvalid             ),
/*  input          */   .S01_AXI_RREADY                  (s01_inf.axi_rready             ),

/*  output         */   .S02_AXI_ARESET_OUT_N            (S02_AXI_ARESET_OUT_N       ),
/*  input          */   .S02_AXI_ACLK                    (s02_inf.axi_aclk           ),
/*  input [0:0]    */   .S02_AXI_AWID                    (s02_inf.axi_awid           ),
/*  input [28:0]   */   .S02_AXI_AWADDR                  (s02_inf.axi_awaddr         ),
/*  input [7:0]    */   .S02_AXI_AWLEN                   (s02_inf.axi_awlen          ),
/*  input [2:0]    */   .S02_AXI_AWSIZE                  (s02_inf.axi_awsize         ),
/*  input [1:0]    */   .S02_AXI_AWBURST                 (s02_inf.axi_awburst        ),
/*  input          */   .S02_AXI_AWLOCK                  (s02_inf.axi_awlock         ),
/*  input [3:0]    */   .S02_AXI_AWCACHE                 (s02_inf.axi_awcache        ),
/*  input [2:0]    */   .S02_AXI_AWPROT                  (s02_inf.axi_awprot         ),
/*  input [3:0]    */   .S02_AXI_AWQOS                   (s02_inf.axi_awqos          ),
/*  input          */   .S02_AXI_AWVALID                 (s02_inf.axi_awvalid        ),
/*  output         */   .S02_AXI_AWREADY                 (s02_inf.axi_awready        ),
/*  input [511:0]  */   .S02_AXI_WDATA                   (s02_inf.axi_wdata          ),
/*  input [63:0]   */   .S02_AXI_WSTRB                   (s02_inf.axi_wstrb          ),
/*  input          */   .S02_AXI_WLAST                   (s02_inf.axi_wlast          ),
/*  input          */   .S02_AXI_WVALID                  (s02_inf.axi_wvalid         ),
/*  output         */   .S02_AXI_WREADY                  (s02_inf.axi_wready         ),
/*  output [0:0]   */   .S02_AXI_BID                     (s02_inf.axi_bid            ),
/*  output [1:0]   */   .S02_AXI_BRESP                   (s02_inf.axi_bresp          ),
/*  output         */   .S02_AXI_BVALID                  (s02_inf.axi_bvalid         ),
/*  input          */   .S02_AXI_BREADY                  (s02_inf.axi_bready         ),
/*  input [0:0]    */   .S02_AXI_ARID                    (s02_inf.axi_arid           ),
/*  input [28:0]   */   .S02_AXI_ARADDR                  (s02_inf.axi_araddr         ),
/*  input [7:0]    */   .S02_AXI_ARLEN                   (s02_inf.axi_arlen          ),
/*  input [2:0]    */   .S02_AXI_ARSIZE                  (s02_inf.axi_arsize         ),
/*  input [1:0]    */   .S02_AXI_ARBURST                 (s02_inf.axi_arburst        ),
/*  input          */   .S02_AXI_ARLOCK                  (s02_inf.axi_arlock         ),
/*  input [3:0]    */   .S02_AXI_ARCACHE                 (s02_inf.axi_arcache        ),
/*  input [2:0]    */   .S02_AXI_ARPROT                  (s02_inf.axi_arprot         ),
/*  input [3:0]    */   .S02_AXI_ARQOS                   (s02_inf.axi_arqos          ),
/*  input          */   .S02_AXI_ARVALID                 (s02_inf.axi_arvalid        ),
/*  output         */   .S02_AXI_ARREADY                 (s02_inf.axi_arready        ),
/*  output [0:0]   */   .S02_AXI_RID                     (s02_inf.axi_rid            ),
/*  output [511:0] */   .S02_AXI_RDATA                   (s02_inf.axi_rdata          ),
/*  output [1:0]   */   .S02_AXI_RRESP                   (s02_inf.axi_rresp          ),
/*  output         */   .S02_AXI_RLAST                   (s02_inf.axi_rlast          ),
/*  output         */   .S02_AXI_RVALID                  (s02_inf.axi_rvalid         ),
/*  input          */   .S02_AXI_RREADY                  (s02_inf.axi_rready         ),
/*  output S01_AXI_*/   .S03_AXI_ARESET_OUT_N            (S03_AXI_ARESET_OUT_N       ),
/*  input          */   .S03_AXI_ACLK                    (s03_inf.axi_aclk               ),
/*  input [0:0]    */   .S03_AXI_AWID                    (s03_inf.axi_awid               ),
/*  input [28:0]   */   .S03_AXI_AWADDR                  (s03_inf.axi_awaddr             ),
/*  input [7:0]    */   .S03_AXI_AWLEN                   (s03_inf.axi_awlen              ),
/*  input [2:0]    */   .S03_AXI_AWSIZE                  (s03_inf.axi_awsize             ),
/*  input [1:0]    */   .S03_AXI_AWBURST                 (s03_inf.axi_awburst            ),
/*  input          */   .S03_AXI_AWLOCK                  (s03_inf.axi_awlock             ),
/*  input [3:0]    */   .S03_AXI_AWCACHE                 (s03_inf.axi_awcache            ),
/*  input [2:0]    */   .S03_AXI_AWPROT                  (s03_inf.axi_awprot             ),
/*  input [3:0]    */   .S03_AXI_AWQOS                   (s03_inf.axi_awqos              ),
/*  input          */   .S03_AXI_AWVALID                 (s03_inf.axi_awvalid            ),
/*  output         */   .S03_AXI_AWREADY                 (s03_inf.axi_awready            ),
/*  input [511:0]  */   .S03_AXI_WDATA                   (s03_inf.axi_wdata              ),
/*  input [63:0]   */   .S03_AXI_WSTRB                   (s03_inf.axi_wstrb              ),
/*  input          */   .S03_AXI_WLAST                   (s03_inf.axi_wlast              ),
/*  input          */   .S03_AXI_WVALID                  (s03_inf.axi_wvalid             ),
/*  output         */   .S03_AXI_WREADY                  (s03_inf.axi_wready             ),
/*  output [0:0]   */   .S03_AXI_BID                     (s03_inf.axi_bid                ),
/*  output [1:0]   */   .S03_AXI_BRESP                   (s03_inf.axi_bresp              ),
/*  output         */   .S03_AXI_BVALID                  (s03_inf.axi_bvalid             ),
/*  input          */   .S03_AXI_BREADY                  (s03_inf.axi_bready             ),
/*  input [0:0]    */   .S03_AXI_ARID                    (s03_inf.axi_arid               ),
/*  input [28:0]   */   .S03_AXI_ARADDR                  (s03_inf.axi_araddr             ),
/*  input [7:0]    */   .S03_AXI_ARLEN                   (s03_inf.axi_arlen              ),
/*  input [2:0]    */   .S03_AXI_ARSIZE                  (s03_inf.axi_arsize             ),
/*  input [1:0]    */   .S03_AXI_ARBURST                 (s03_inf.axi_arburst            ),
/*  input          */   .S03_AXI_ARLOCK                  (s03_inf.axi_arlock             ),
/*  input [3:0]    */   .S03_AXI_ARCACHE                 (s03_inf.axi_arcache            ),
/*  input [2:0]    */   .S03_AXI_ARPROT                  (s03_inf.axi_arprot             ),
/*  input [3:0]    */   .S03_AXI_ARQOS                   (s03_inf.axi_arqos              ),
/*  input          */   .S03_AXI_ARVALID                 (s03_inf.axi_arvalid            ),
/*  output         */   .S03_AXI_ARREADY                 (s03_inf.axi_arready            ),
/*  output [0:0]   */   .S03_AXI_RID                     (s03_inf.axi_rid                ),
/*  output [511:0] */   .S03_AXI_RDATA                   (s03_inf.axi_rdata              ),
/*  output [1:0]   */   .S03_AXI_RRESP                   (s03_inf.axi_rresp              ),
/*  output         */   .S03_AXI_RLAST                   (s03_inf.axi_rlast              ),
/*  output         */   .S03_AXI_RVALID                  (s03_inf.axi_rvalid             ),
/*  input          */   .S03_AXI_RREADY                  (s03_inf.axi_rready             ),

/*  output         */   .S04_AXI_ARESET_OUT_N            (S04_AXI_ARESET_OUT_N       ),
/*  input          */   .S04_AXI_ACLK                    (s04_inf.axi_aclk           ),
/*  input [0:0]    */   .S04_AXI_AWID                    (s04_inf.axi_awid           ),
/*  input [28:0]   */   .S04_AXI_AWADDR                  (s04_inf.axi_awaddr         ),
/*  input [7:0]    */   .S04_AXI_AWLEN                   (s04_inf.axi_awlen          ),
/*  input [2:0]    */   .S04_AXI_AWSIZE                  (s04_inf.axi_awsize         ),
/*  input [1:0]    */   .S04_AXI_AWBURST                 (s04_inf.axi_awburst        ),
/*  input          */   .S04_AXI_AWLOCK                  (s04_inf.axi_awlock         ),
/*  input [3:0]    */   .S04_AXI_AWCACHE                 (s04_inf.axi_awcache        ),
/*  input [2:0]    */   .S04_AXI_AWPROT                  (s04_inf.axi_awprot         ),
/*  input [3:0]    */   .S04_AXI_AWQOS                   (s04_inf.axi_awqos          ),
/*  input          */   .S04_AXI_AWVALID                 (s04_inf.axi_awvalid        ),
/*  output         */   .S04_AXI_AWREADY                 (s04_inf.axi_awready        ),
/*  input [511:0]  */   .S04_AXI_WDATA                   (s04_inf.axi_wdata          ),
/*  input [63:0]   */   .S04_AXI_WSTRB                   (s04_inf.axi_wstrb          ),
/*  input          */   .S04_AXI_WLAST                   (s04_inf.axi_wlast          ),
/*  input          */   .S04_AXI_WVALID                  (s04_inf.axi_wvalid         ),
/*  output         */   .S04_AXI_WREADY                  (s04_inf.axi_wready         ),
/*  output [0:0]   */   .S04_AXI_BID                     (s04_inf.axi_bid            ),
/*  output [1:0]   */   .S04_AXI_BRESP                   (s04_inf.axi_bresp          ),
/*  output         */   .S04_AXI_BVALID                  (s04_inf.axi_bvalid         ),
/*  input          */   .S04_AXI_BREADY                  (s04_inf.axi_bready         ),
/*  input [0:0]    */   .S04_AXI_ARID                    (s04_inf.axi_arid           ),
/*  input [28:0]   */   .S04_AXI_ARADDR                  (s04_inf.axi_araddr         ),
/*  input [7:0]    */   .S04_AXI_ARLEN                   (s04_inf.axi_arlen          ),
/*  input [2:0]    */   .S04_AXI_ARSIZE                  (s04_inf.axi_arsize         ),
/*  input [1:0]    */   .S04_AXI_ARBURST                 (s04_inf.axi_arburst        ),
/*  input          */   .S04_AXI_ARLOCK                  (s04_inf.axi_arlock         ),
/*  input [3:0]    */   .S04_AXI_ARCACHE                 (s04_inf.axi_arcache        ),
/*  input [2:0]    */   .S04_AXI_ARPROT                  (s04_inf.axi_arprot         ),
/*  input [3:0]    */   .S04_AXI_ARQOS                   (s04_inf.axi_arqos          ),
/*  input          */   .S04_AXI_ARVALID                 (s04_inf.axi_arvalid        ),
/*  output         */   .S04_AXI_ARREADY                 (s04_inf.axi_arready        ),
/*  output [0:0]   */   .S04_AXI_RID                     (s04_inf.axi_rid            ),
/*  output [511:0] */   .S04_AXI_RDATA                   (s04_inf.axi_rdata          ),
/*  output [1:0]   */   .S04_AXI_RRESP                   (s04_inf.axi_rresp          ),
/*  output         */   .S04_AXI_RLAST                   (s04_inf.axi_rlast          ),
/*  output         */   .S04_AXI_RVALID                  (s04_inf.axi_rvalid         ),
/*  input          */   .S04_AXI_RREADY                  (s04_inf.axi_rready         ),
/*  output S01_AXI_*/   .S05_AXI_ARESET_OUT_N            (S05_AXI_ARESET_OUT_N       ),
/*  input          */   .S05_AXI_ACLK                    (s05_inf.axi_aclk               ),
/*  input [0:0]    */   .S05_AXI_AWID                    (s05_inf.axi_awid               ),
/*  input [28:0]   */   .S05_AXI_AWADDR                  (s05_inf.axi_awaddr             ),
/*  input [7:0]    */   .S05_AXI_AWLEN                   (s05_inf.axi_awlen              ),
/*  input [2:0]    */   .S05_AXI_AWSIZE                  (s05_inf.axi_awsize             ),
/*  input [1:0]    */   .S05_AXI_AWBURST                 (s05_inf.axi_awburst            ),
/*  input          */   .S05_AXI_AWLOCK                  (s05_inf.axi_awlock             ),
/*  input [3:0]    */   .S05_AXI_AWCACHE                 (s05_inf.axi_awcache            ),
/*  input [2:0]    */   .S05_AXI_AWPROT                  (s05_inf.axi_awprot             ),
/*  input [3:0]    */   .S05_AXI_AWQOS                   (s05_inf.axi_awqos              ),
/*  input          */   .S05_AXI_AWVALID                 (s05_inf.axi_awvalid            ),
/*  output         */   .S05_AXI_AWREADY                 (s05_inf.axi_awready            ),
/*  input [511:0]  */   .S05_AXI_WDATA                   (s05_inf.axi_wdata              ),
/*  input [63:0]   */   .S05_AXI_WSTRB                   (s05_inf.axi_wstrb              ),
/*  input          */   .S05_AXI_WLAST                   (s05_inf.axi_wlast              ),
/*  input          */   .S05_AXI_WVALID                  (s05_inf.axi_wvalid             ),
/*  output         */   .S05_AXI_WREADY                  (s05_inf.axi_wready             ),
/*  output [0:0]   */   .S05_AXI_BID                     (s05_inf.axi_bid                ),
/*  output [1:0]   */   .S05_AXI_BRESP                   (s05_inf.axi_bresp              ),
/*  output         */   .S05_AXI_BVALID                  (s05_inf.axi_bvalid             ),
/*  input          */   .S05_AXI_BREADY                  (s05_inf.axi_bready             ),
/*  input [0:0]    */   .S05_AXI_ARID                    (s05_inf.axi_arid               ),
/*  input [28:0]   */   .S05_AXI_ARADDR                  (s05_inf.axi_araddr             ),
/*  input [7:0]    */   .S05_AXI_ARLEN                   (s05_inf.axi_arlen              ),
/*  input [2:0]    */   .S05_AXI_ARSIZE                  (s05_inf.axi_arsize             ),
/*  input [1:0]    */   .S05_AXI_ARBURST                 (s05_inf.axi_arburst            ),
/*  input          */   .S05_AXI_ARLOCK                  (s05_inf.axi_arlock             ),
/*  input [3:0]    */   .S05_AXI_ARCACHE                 (s05_inf.axi_arcache            ),
/*  input [2:0]    */   .S05_AXI_ARPROT                  (s05_inf.axi_arprot             ),
/*  input [3:0]    */   .S05_AXI_ARQOS                   (s05_inf.axi_arqos              ),
/*  input          */   .S05_AXI_ARVALID                 (s05_inf.axi_arvalid            ),
/*  output         */   .S05_AXI_ARREADY                 (s05_inf.axi_arready            ),
/*  output [0:0]   */   .S05_AXI_RID                     (s05_inf.axi_rid                ),
/*  output [511:0] */   .S05_AXI_RDATA                   (s05_inf.axi_rdata              ),
/*  output [1:0]   */   .S05_AXI_RRESP                   (s05_inf.axi_rresp              ),
/*  output         */   .S05_AXI_RLAST                   (s05_inf.axi_rlast              ),
/*  output         */   .S05_AXI_RVALID                  (s05_inf.axi_rvalid             ),
/*  input          */   .S05_AXI_RREADY                  (s05_inf.axi_rready             ),

/*  output         */   .S06_AXI_ARESET_OUT_N            (S06_AXI_ARESET_OUT_N       ),
/*  input          */   .S06_AXI_ACLK                    (s06_inf.axi_aclk           ),
/*  input [0:0]    */   .S06_AXI_AWID                    (s06_inf.axi_awid           ),
/*  input [28:0]   */   .S06_AXI_AWADDR                  (s06_inf.axi_awaddr         ),
/*  input [7:0]    */   .S06_AXI_AWLEN                   (s06_inf.axi_awlen          ),
/*  input [2:0]    */   .S06_AXI_AWSIZE                  (s06_inf.axi_awsize         ),
/*  input [1:0]    */   .S06_AXI_AWBURST                 (s06_inf.axi_awburst        ),
/*  input          */   .S06_AXI_AWLOCK                  (s06_inf.axi_awlock         ),
/*  input [3:0]    */   .S06_AXI_AWCACHE                 (s06_inf.axi_awcache        ),
/*  input [2:0]    */   .S06_AXI_AWPROT                  (s06_inf.axi_awprot         ),
/*  input [3:0]    */   .S06_AXI_AWQOS                   (s06_inf.axi_awqos          ),
/*  input          */   .S06_AXI_AWVALID                 (s06_inf.axi_awvalid        ),
/*  output         */   .S06_AXI_AWREADY                 (s06_inf.axi_awready        ),
/*  input [511:0]  */   .S06_AXI_WDATA                   (s06_inf.axi_wdata          ),
/*  input [63:0]   */   .S06_AXI_WSTRB                   (s06_inf.axi_wstrb          ),
/*  input          */   .S06_AXI_WLAST                   (s06_inf.axi_wlast          ),
/*  input          */   .S06_AXI_WVALID                  (s06_inf.axi_wvalid         ),
/*  output         */   .S06_AXI_WREADY                  (s06_inf.axi_wready         ),
/*  output [0:0]   */   .S06_AXI_BID                     (s06_inf.axi_bid            ),
/*  output [1:0]   */   .S06_AXI_BRESP                   (s06_inf.axi_bresp          ),
/*  output         */   .S06_AXI_BVALID                  (s06_inf.axi_bvalid         ),
/*  input          */   .S06_AXI_BREADY                  (s06_inf.axi_bready         ),
/*  input [0:0]    */   .S06_AXI_ARID                    (s06_inf.axi_arid           ),
/*  input [28:0]   */   .S06_AXI_ARADDR                  (s06_inf.axi_araddr         ),
/*  input [7:0]    */   .S06_AXI_ARLEN                   (s06_inf.axi_arlen          ),
/*  input [2:0]    */   .S06_AXI_ARSIZE                  (s06_inf.axi_arsize         ),
/*  input [1:0]    */   .S06_AXI_ARBURST                 (s06_inf.axi_arburst        ),
/*  input          */   .S06_AXI_ARLOCK                  (s06_inf.axi_arlock         ),
/*  input [3:0]    */   .S06_AXI_ARCACHE                 (s06_inf.axi_arcache        ),
/*  input [2:0]    */   .S06_AXI_ARPROT                  (s06_inf.axi_arprot         ),
/*  input [3:0]    */   .S06_AXI_ARQOS                   (s06_inf.axi_arqos          ),
/*  input          */   .S06_AXI_ARVALID                 (s06_inf.axi_arvalid        ),
/*  output         */   .S06_AXI_ARREADY                 (s06_inf.axi_arready        ),
/*  output [0:0]   */   .S06_AXI_RID                     (s06_inf.axi_rid            ),
/*  output [511:0] */   .S06_AXI_RDATA                   (s06_inf.axi_rdata          ),
/*  output [1:0]   */   .S06_AXI_RRESP                   (s06_inf.axi_rresp          ),
/*  output         */   .S06_AXI_RLAST                   (s06_inf.axi_rlast          ),
/*  output         */   .S06_AXI_RVALID                  (s06_inf.axi_rvalid         ),
/*  input          */   .S06_AXI_RREADY                  (s06_inf.axi_rready         ),
/*  output S01_AXI_*/   .S07_AXI_ARESET_OUT_N            (S07_AXI_ARESET_OUT_N       ),
/*  input          */   .S07_AXI_ACLK                    (s07_inf.axi_aclk               ),
/*  input [0:0]    */   .S07_AXI_AWID                    (s07_inf.axi_awid               ),
/*  input [28:0]   */   .S07_AXI_AWADDR                  (s07_inf.axi_awaddr             ),
/*  input [7:0]    */   .S07_AXI_AWLEN                   (s07_inf.axi_awlen              ),
/*  input [2:0]    */   .S07_AXI_AWSIZE                  (s07_inf.axi_awsize             ),
/*  input [1:0]    */   .S07_AXI_AWBURST                 (s07_inf.axi_awburst            ),
/*  input          */   .S07_AXI_AWLOCK                  (s07_inf.axi_awlock             ),
/*  input [3:0]    */   .S07_AXI_AWCACHE                 (s07_inf.axi_awcache            ),
/*  input [2:0]    */   .S07_AXI_AWPROT                  (s07_inf.axi_awprot             ),
/*  input [3:0]    */   .S07_AXI_AWQOS                   (s07_inf.axi_awqos              ),
/*  input          */   .S07_AXI_AWVALID                 (s07_inf.axi_awvalid            ),
/*  output         */   .S07_AXI_AWREADY                 (s07_inf.axi_awready            ),
/*  input [511:0]  */   .S07_AXI_WDATA                   (s07_inf.axi_wdata              ),
/*  input [63:0]   */   .S07_AXI_WSTRB                   (s07_inf.axi_wstrb              ),
/*  input          */   .S07_AXI_WLAST                   (s07_inf.axi_wlast              ),
/*  input          */   .S07_AXI_WVALID                  (s07_inf.axi_wvalid             ),
/*  output         */   .S07_AXI_WREADY                  (s07_inf.axi_wready             ),
/*  output [0:0]   */   .S07_AXI_BID                     (s07_inf.axi_bid                ),
/*  output [1:0]   */   .S07_AXI_BRESP                   (s07_inf.axi_bresp              ),
/*  output         */   .S07_AXI_BVALID                  (s07_inf.axi_bvalid             ),
/*  input          */   .S07_AXI_BREADY                  (s07_inf.axi_bready             ),
/*  input [0:0]    */   .S07_AXI_ARID                    (s07_inf.axi_arid               ),
/*  input [28:0]   */   .S07_AXI_ARADDR                  (s07_inf.axi_araddr             ),
/*  input [7:0]    */   .S07_AXI_ARLEN                   (s07_inf.axi_arlen              ),
/*  input [2:0]    */   .S07_AXI_ARSIZE                  (s07_inf.axi_arsize             ),
/*  input [1:0]    */   .S07_AXI_ARBURST                 (s07_inf.axi_arburst            ),
/*  input          */   .S07_AXI_ARLOCK                  (s07_inf.axi_arlock             ),
/*  input [3:0]    */   .S07_AXI_ARCACHE                 (s07_inf.axi_arcache            ),
/*  input [2:0]    */   .S07_AXI_ARPROT                  (s07_inf.axi_arprot             ),
/*  input [3:0]    */   .S07_AXI_ARQOS                   (s07_inf.axi_arqos              ),
/*  input          */   .S07_AXI_ARVALID                 (s07_inf.axi_arvalid            ),
/*  output         */   .S07_AXI_ARREADY                 (s07_inf.axi_arready            ),
/*  output [0:0]   */   .S07_AXI_RID                     (s07_inf.axi_rid                ),
/*  output [511:0] */   .S07_AXI_RDATA                   (s07_inf.axi_rdata              ),
/*  output [1:0]   */   .S07_AXI_RRESP                   (s07_inf.axi_rresp              ),
/*  output         */   .S07_AXI_RLAST                   (s07_inf.axi_rlast              ),
/*  output         */   .S07_AXI_RVALID                  (s07_inf.axi_rvalid             ),
/*  input          */   .S07_AXI_RREADY                  (s07_inf.axi_rready             ),


/*  output         */   .M00_AXI_ARESET_OUT_N            (M00_AXI_ARESET_OUT_N           ),
/*  input          */   .M00_AXI_ACLK                    (m00_inf.axi_aclk               ),
/*  output [3:0]   */   .M00_AXI_AWID                    (m00_inf.axi_awid               ),
/*  output [28:0]  */   .M00_AXI_AWADDR                  (m00_inf.axi_awaddr             ),
/*  output [7:0]   */   .M00_AXI_AWLEN                   (m00_inf.axi_awlen              ),
/*  output [2:0]   */   .M00_AXI_AWSIZE                  (m00_inf.axi_awsize             ),
/*  output [1:0]   */   .M00_AXI_AWBURST                 (m00_inf.axi_awburst            ),
/*  output         */   .M00_AXI_AWLOCK                  (m00_inf.axi_awlock             ),
/*  output [3:0]   */   .M00_AXI_AWCACHE                 (m00_inf.axi_awcache            ),
/*  output [2:0]   */   .M00_AXI_AWPROT                  (m00_inf.axi_awprot             ),
/*  output [3:0]   */   .M00_AXI_AWQOS                   (m00_inf.axi_awqos              ),
/*  output         */   .M00_AXI_AWVALID                 (m00_inf.axi_awvalid            ),
/*  input          */   .M00_AXI_AWREADY                 (m00_inf.axi_awready            ),
/*  output [511:0] */   .M00_AXI_WDATA                   (m00_inf.axi_wdata              ),
/*  output [63:0]  */   .M00_AXI_WSTRB                   (m00_inf.axi_wstrb              ),
/*  output         */   .M00_AXI_WLAST                   (m00_inf.axi_wlast              ),
/*  output         */   .M00_AXI_WVALID                  (m00_inf.axi_wvalid             ),
/*  input          */   .M00_AXI_WREADY                  (m00_inf.axi_wready             ),
/*  input [3:0]    */   .M00_AXI_BID                     (m00_inf.axi_bid                ),
/*  input [1:0]    */   .M00_AXI_BRESP                   (m00_inf.axi_bresp              ),
/*  input          */   .M00_AXI_BVALID                  (m00_inf.axi_bvalid             ),
/*  output         */   .M00_AXI_BREADY                  (m00_inf.axi_bready             ),
/*  output [3:0]   */   .M00_AXI_ARID                    (m00_inf.axi_arid               ),
/*  output [28:0]  */   .M00_AXI_ARADDR                  (m00_inf.axi_araddr             ),
/*  output [7:0]   */   .M00_AXI_ARLEN                   (m00_inf.axi_arlen              ),
/*  output [2:0]   */   .M00_AXI_ARSIZE                  (m00_inf.axi_arsize             ),
/*  output [1:0]   */   .M00_AXI_ARBURST                 (m00_inf.axi_arburst            ),
/*  output         */   .M00_AXI_ARLOCK                  (m00_inf.axi_arlock             ),
/*  output [3:0]   */   .M00_AXI_ARCACHE                 (m00_inf.axi_arcache            ),
/*  output [2:0]   */   .M00_AXI_ARPROT                  (m00_inf.axi_arprot             ),
/*  output [3:0]   */   .M00_AXI_ARQOS                   (m00_inf.axi_arqos              ),
/*  output         */   .M00_AXI_ARVALID                 (m00_inf.axi_arvalid            ),
/*  input          */   .M00_AXI_ARREADY                 (m00_inf.axi_arready            ),
/*  input [3:0]    */   .M00_AXI_RID                     (m00_inf.axi_rid                ),
/*  input [511:0]  */   .M00_AXI_RDATA                   (m00_inf.axi_rdata              ),
/*  input [1:0]    */   .M00_AXI_RRESP                   (m00_inf.axi_rresp              ),
/*  input          */   .M00_AXI_RLAST                   (m00_inf.axi_rlast              ),
/*  input          */   .M00_AXI_RVALID                  (m00_inf.axi_rvalid             ),
/*  output         */   .M00_AXI_RREADY                  (m00_inf.axi_rready             )
);
end
endgenerate

assign s00_inf.axi_wevld   = m00_inf.axi_wevld    ;
assign s00_inf.axi_weresp  = m00_inf.axi_weresp   ;
assign s00_inf.axi_revld   = m00_inf.axi_revld    ;
assign s00_inf.axi_reresp  = m00_inf.axi_reresp   ;

assign s01_inf.axi_wevld   = m00_inf.axi_wevld    ;
assign s01_inf.axi_weresp  = m00_inf.axi_weresp   ;
assign s01_inf.axi_revld   = m00_inf.axi_revld    ;
assign s01_inf.axi_reresp  = m00_inf.axi_reresp   ;

assign s02_inf.axi_wevld   = m00_inf.axi_wevld    ;
assign s02_inf.axi_weresp  = m00_inf.axi_weresp   ;
assign s02_inf.axi_revld   = m00_inf.axi_revld    ;
assign s02_inf.axi_reresp  = m00_inf.axi_reresp   ;

assign s03_inf.axi_wevld   = m00_inf.axi_wevld    ;
assign s03_inf.axi_weresp  = m00_inf.axi_weresp   ;
assign s03_inf.axi_revld   = m00_inf.axi_revld    ;
assign s03_inf.axi_reresp  = m00_inf.axi_reresp   ;

assign s04_inf.axi_wevld   = m00_inf.axi_wevld    ;
assign s04_inf.axi_weresp  = m00_inf.axi_weresp   ;
assign s04_inf.axi_revld   = m00_inf.axi_revld    ;
assign s04_inf.axi_reresp  = m00_inf.axi_reresp   ;

assign s05_inf.axi_wevld   = m00_inf.axi_wevld    ;
assign s05_inf.axi_weresp  = m00_inf.axi_weresp   ;
assign s05_inf.axi_revld   = m00_inf.axi_revld    ;
assign s05_inf.axi_reresp  = m00_inf.axi_reresp   ;

assign s06_inf.axi_wevld   = m00_inf.axi_wevld    ;
assign s06_inf.axi_weresp  = m00_inf.axi_weresp   ;
assign s06_inf.axi_revld   = m00_inf.axi_revld    ;
assign s06_inf.axi_reresp  = m00_inf.axi_reresp   ;

assign s07_inf.axi_wevld   = m00_inf.axi_wevld    ;
assign s07_inf.axi_weresp  = m00_inf.axi_weresp   ;
assign s07_inf.axi_revld   = m00_inf.axi_revld    ;
assign s07_inf.axi_reresp  = m00_inf.axi_reresp   ;

endmodule
