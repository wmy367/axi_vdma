/**********************************************
______________                ______________
______________ \  /\  /|\  /| ______________
______________  \/  \/ | \/ | ______________
descript:
    axi4 write read lock ,pend each other
author : Young
Version: VERA.0.0
creaded: 2016/8/29 下午3:29:24
madified:
***********************************************/
`timescale 1ns/1ps
module axi4_interconnect_wrap (
    input          INTERCONNECT_ACLK    ,
    input          INTERCONNECT_ARESETN ,
    output         S00_AXI_ARESET_OUT_N ,
    output         S01_AXI_ARESET_OUT_N ,
    output         M00_AXI_ARESET_OUT_N ,
    axi_inf.slaver s00_inf  ,
    axi_inf.slaver s01_inf  ,
    axi_inf.master m00_inf
);

AXI4_INFCNT AXI4_INFCNT_inst(
/*  input          */   .INTERCONNECT_ACLK               (INTERCONNECT_ACLK          ),
/*  input          */   .INTERCONNECT_ARESETN            (INTERCONNECT_ARESETN       ),
/*  output         */   .S00_AXI_ARESET_OUT_N            (S00_AXI_ARESET_OUT_N       ),
/*  input          */   .S00_AXI_ACLK                    (s00_inf.axi_aclk           ),
/*  input [0:0]    */   .S00_AXI_AWID                    (s00_inf.axi_awid           ),
/*  input [28:0]   */   .S00_AXI_AWADDR                  (s00_inf.axi_awaddr         ),
/*  input [7:0]    */   .S00_AXI_AWLEN                   (s00_inf.axi_awlen          ),
/*  input [2:0]    */   .S00_AXI_AWSIZE                  (s00_inf.axi_awsize         ),
/*  input [1:0]    */   .S00_AXI_AWBURST                 (s00_inf.axi_awburst        ),
/*  input          */   .S00_AXI_AWLOCK                  (s00_inf.axi_awlock         ),
/*  input [3:0]    */   .S00_AXI_AWCACHE                 (s00_inf.axi_awcache        ),
/*  input [2:0]    */   .S00_AXI_AWPROT                  (s00_inf.axi_awprot         ),
/*  input [3:0]    */   .S00_AXI_AWQOS                   (s00_inf.axi_awqos          ),
/*  input          */   .S00_AXI_AWVALID                 (s00_inf.axi_awvalid        ),
/*  output         */   .S00_AXI_AWREADY                 (s00_inf.axi_awready        ),
/*  input [255:0]  */   .S00_AXI_WDATA                   (s00_inf.axi_wdata          ),
/*  input [31:0]   */   .S00_AXI_WSTRB                   (s00_inf.axi_wstrb          ),
/*  input          */   .S00_AXI_WLAST                   (s00_inf.axi_wlast          ),
/*  input          */   .S00_AXI_WVALID                  (s00_inf.axi_wvalid         ),
/*  output         */   .S00_AXI_WREADY                  (s00_inf.axi_wready         ),
/*  output [0:0]   */   .S00_AXI_BID                     (s00_inf.axi_bid            ),
/*  output [1:0]   */   .S00_AXI_BRESP                   (s00_inf.axi_bresp          ),
/*  output         */   .S00_AXI_BVALID                  (s00_inf.axi_bvalid         ),
/*  input          */   .S00_AXI_BREADY                  (s00_inf.axi_bready         ),
/*  input [0:0]    */   .S00_AXI_ARID                    (s00_inf.axi_arid           ),
/*  input [28:0]   */   .S00_AXI_ARADDR                  (s00_inf.axi_araddr         ),
/*  input [7:0]    */   .S00_AXI_ARLEN                   (s00_inf.axi_arlen          ),
/*  input [2:0]    */   .S00_AXI_ARSIZE                  (s00_inf.axi_arsize         ),
/*  input [1:0]    */   .S00_AXI_ARBURST                 (s00_inf.axi_arburst        ),
/*  input          */   .S00_AXI_ARLOCK                  (s00_inf.axi_arlock         ),
/*  input [3:0]    */   .S00_AXI_ARCACHE                 (s00_inf.axi_arcache        ),
/*  input [2:0]    */   .S00_AXI_ARPROT                  (s00_inf.axi_arprot         ),
/*  input [3:0]    */   .S00_AXI_ARQOS                   (s00_inf.axi_arqos          ),
/*  input          */   .S00_AXI_ARVALID                 (s00_inf.axi_arvalid        ),
/*  output         */   .S00_AXI_ARREADY                 (s00_inf.axi_arready        ),
/*  output [0:0]   */   .S00_AXI_RID                     (s00_inf.axi_rid            ),
/*  output [255:0] */   .S00_AXI_RDATA                   (s00_inf.axi_rdata          ),
/*  output [1:0]   */   .S00_AXI_RRESP                   (s00_inf.axi_rresp          ),
/*  output         */   .S00_AXI_RLAST                   (s00_inf.axi_rlast          ),
/*  output         */   .S00_AXI_RVALID                  (s00_inf.axi_rvalid         ),
/*  input          */   .S00_AXI_RREADY                  (s00_inf.axi_rready         ),
/*  output S01_AXI_*/   .S01_AXI_ARESET_OUT_N            (S01_AXI_ARESET_OUT_N       ),
/*  input          */   .S01_AXI_ACLK                    (s01_inf.axi_aclk               ),
/*  input [0:0]    */   .S01_AXI_AWID                    (s01_inf.axi_awid               ),
/*  input [28:0]   */   .S01_AXI_AWADDR                  (s01_inf.axi_awaddr             ),
/*  input [7:0]    */   .S01_AXI_AWLEN                   (s01_inf.axi_awlen              ),
/*  input [2:0]    */   .S01_AXI_AWSIZE                  (s01_inf.axi_awsize             ),
/*  input [1:0]    */   .S01_AXI_AWBURST                 (s01_inf.axi_awburst            ),
/*  input          */   .S01_AXI_AWLOCK                  (s01_inf.axi_awlock             ),
/*  input [3:0]    */   .S01_AXI_AWCACHE                 (s01_inf.axi_awcache            ),
/*  input [2:0]    */   .S01_AXI_AWPROT                  (s01_inf.axi_awprot             ),
/*  input [3:0]    */   .S01_AXI_AWQOS                   (s01_inf.axi_awqos              ),
/*  input          */   .S01_AXI_AWVALID                 (s01_inf.axi_awvalid            ),
/*  output         */   .S01_AXI_AWREADY                 (s01_inf.axi_awready            ),
/*  input [255:0]  */   .S01_AXI_WDATA                   (s01_inf.axi_wdata              ),
/*  input [31:0]   */   .S01_AXI_WSTRB                   (s01_inf.axi_wstrb              ),
/*  input          */   .S01_AXI_WLAST                   (s01_inf.axi_wlast              ),
/*  input          */   .S01_AXI_WVALID                  (s01_inf.axi_wvalid             ),
/*  output         */   .S01_AXI_WREADY                  (s01_inf.axi_wready             ),
/*  output [0:0]   */   .S01_AXI_BID                     (s01_inf.axi_bid                ),
/*  output [1:0]   */   .S01_AXI_BRESP                   (s01_inf.axi_bresp              ),
/*  output         */   .S01_AXI_BVALID                  (s01_inf.axi_bvalid             ),
/*  input          */   .S01_AXI_BREADY                  (s01_inf.axi_bready             ),
/*  input [0:0]    */   .S01_AXI_ARID                    (s01_inf.axi_arid               ),
/*  input [28:0]   */   .S01_AXI_ARADDR                  (s01_inf.axi_araddr             ),
/*  input [7:0]    */   .S01_AXI_ARLEN                   (s01_inf.axi_arlen              ),
/*  input [2:0]    */   .S01_AXI_ARSIZE                  (s01_inf.axi_arsize             ),
/*  input [1:0]    */   .S01_AXI_ARBURST                 (s01_inf.axi_arburst            ),
/*  input          */   .S01_AXI_ARLOCK                  (s01_inf.axi_arlock             ),
/*  input [3:0]    */   .S01_AXI_ARCACHE                 (s01_inf.axi_arcache            ),
/*  input [2:0]    */   .S01_AXI_ARPROT                  (s01_inf.axi_arprot             ),
/*  input [3:0]    */   .S01_AXI_ARQOS                   (s01_inf.axi_arqos              ),
/*  input          */   .S01_AXI_ARVALID                 (s01_inf.axi_arvalid            ),
/*  output         */   .S01_AXI_ARREADY                 (s01_inf.axi_arready            ),
/*  output [0:0]   */   .S01_AXI_RID                     (s01_inf.axi_rid                ),
/*  output [255:0] */   .S01_AXI_RDATA                   (s01_inf.axi_rdata              ),
/*  output [1:0]   */   .S01_AXI_RRESP                   (s01_inf.axi_rresp              ),
/*  output         */   .S01_AXI_RLAST                   (s01_inf.axi_rlast              ),
/*  output         */   .S01_AXI_RVALID                  (s01_inf.axi_rvalid             ),
/*  input          */   .S01_AXI_RREADY                  (s01_inf.axi_rready             ),
/*  output         */   .M00_AXI_ARESET_OUT_N            (M00_AXI_ARESET_OUT_N           ),
/*  input          */   .M00_AXI_ACLK                    (m00_inf.axi_aclk               ),
/*  output [3:0]   */   .M00_AXI_AWID                    (m00_inf.axi_awid               ),
/*  output [28:0]  */   .M00_AXI_AWADDR                  (m00_inf.axi_awaddr             ),
/*  output [7:0]   */   .M00_AXI_AWLEN                   (m00_inf.axi_awlen              ),
/*  output [2:0]   */   .M00_AXI_AWSIZE                  (m00_inf.axi_awsize             ),
/*  output [1:0]   */   .M00_AXI_AWBURST                 (m00_inf.axi_awburst            ),
/*  output         */   .M00_AXI_AWLOCK                  (m00_inf.axi_awlock             ),
/*  output [3:0]   */   .M00_AXI_AWCACHE                 (m00_inf.axi_awcache            ),
/*  output [2:0]   */   .M00_AXI_AWPROT                  (m00_inf.axi_awprot             ),
/*  output [3:0]   */   .M00_AXI_AWQOS                   (m00_inf.axi_awqos              ),
/*  output         */   .M00_AXI_AWVALID                 (m00_inf.axi_awvalid            ),
/*  input          */   .M00_AXI_AWREADY                 (m00_inf.axi_awready            ),
/*  output [255:0] */   .M00_AXI_WDATA                   (m00_inf.axi_wdata              ),
/*  output [31:0]  */   .M00_AXI_WSTRB                   (m00_inf.axi_wstrb              ),
/*  output         */   .M00_AXI_WLAST                   (m00_inf.axi_wlast              ),
/*  output         */   .M00_AXI_WVALID                  (m00_inf.axi_wvalid             ),
/*  input          */   .M00_AXI_WREADY                  (m00_inf.axi_wready             ),
/*  input [3:0]    */   .M00_AXI_BID                     (m00_inf.axi_bid                ),
/*  input [1:0]    */   .M00_AXI_BRESP                   (m00_inf.axi_bresp              ),
/*  input          */   .M00_AXI_BVALID                  (m00_inf.axi_bvalid             ),
/*  output         */   .M00_AXI_BREADY                  (m00_inf.axi_bready             ),
/*  output [3:0]   */   .M00_AXI_ARID                    (m00_inf.axi_arid               ),
/*  output [28:0]  */   .M00_AXI_ARADDR                  (m00_inf.axi_araddr             ),
/*  output [7:0]   */   .M00_AXI_ARLEN                   (m00_inf.axi_arlen              ),
/*  output [2:0]   */   .M00_AXI_ARSIZE                  (m00_inf.axi_arsize             ),
/*  output [1:0]   */   .M00_AXI_ARBURST                 (m00_inf.axi_arburst            ),
/*  output         */   .M00_AXI_ARLOCK                  (m00_inf.axi_arlock             ),
/*  output [3:0]   */   .M00_AXI_ARCACHE                 (m00_inf.axi_arcache            ),
/*  output [2:0]   */   .M00_AXI_ARPROT                  (m00_inf.axi_arprot             ),
/*  output [3:0]   */   .M00_AXI_ARQOS                   (m00_inf.axi_arqos              ),
/*  output         */   .M00_AXI_ARVALID                 (m00_inf.axi_arvalid            ),
/*  input          */   .M00_AXI_ARREADY                 (m00_inf.axi_arready            ),
/*  input [3:0]    */   .M00_AXI_RID                     (m00_inf.axi_rid                ),
/*  input [255:0]  */   .M00_AXI_RDATA                   (m00_inf.axi_rdata              ),
/*  input [1:0]    */   .M00_AXI_RRESP                   (m00_inf.axi_rresp              ),
/*  input          */   .M00_AXI_RLAST                   (m00_inf.axi_rlast              ),
/*  input          */   .M00_AXI_RVALID                  (m00_inf.axi_rvalid             ),
/*  output         */   .M00_AXI_RREADY                  (m00_inf.axi_rready             )
);

endmodule
